module ADD(
    input [15:0]x,
    input [15:0]y,
    output [15:0] res
);
assign res = x + y;
endmodule
